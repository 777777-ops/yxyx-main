//二进制4位的7位数码管()
module bcd7seg(
  input  [3:0] b,
  output reg [7:0] h
);
  always @(*) begin
    case(b)
      4'h0: h = ~(8'b11111101);  
      4'h1: h = ~(8'b01100000);  
      4'h2: h = ~(8'b11011010);  
      4'h3: h = ~(8'b11110010); 
      4'h4: h = ~(8'b01100110); 
      4'h5: h = ~(8'b10110110); 
      4'h6: h = ~(8'b10111110); 
      4'h7: h = ~(8'b11100000);
      4'h8: h = ~(8'b11111111);
      /* 
      4'h9: h = 7'b1101111;  
      4'hA: h = 7'b1110111;  
      4'hB: h = 7'b1111100;  
      4'hC: h = 7'b0111001;  
      4'hD: h = 7'b1011110;  
      4'hE: h = 7'b1111001;  
      4'hF: h = 7'b1110001;  
      */
      default: h = 8'b00000010; 
    endcase
  end
endmodule




